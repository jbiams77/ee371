module seg7(num, out);
